`define numPorts 16
